module or_gate
(
	input_1,
	input_2,
	or_result
);

	input input_1;
	input input_2;
	output or_result;

	assign or_result = input_1 | input_2;

endmodule
