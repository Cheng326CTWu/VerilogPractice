module not_gate
(
	input_1,
	not_result
);

	input input_1;
	output not_result;

	assign not_result = !input_1;

endmodule
