module and_gate 
(
    input_1,
    input_2,
    and_result
);

	input  input_1;
  	input  input_2;
  	output and_result;
   
  	assign and_result = input_1 & input_2;
 
endmodule // and_gate
